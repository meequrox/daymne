module handler

pub fn main(help_msg string) {
	println(help_msg)
}
